conectix             ,Txvbox   Wi2k     �      �     ����E$�D�C�zD�*��B                                                                                                                                                                                                                                                                                                                                                                                                                                            cxsparse��������                 ���v                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            conectix             ,Txvbox   Wi2k     �      �     ����E$�D�C�zD�*��B                                                                                                                                                                                                                                                                                                                                                                                                                                            